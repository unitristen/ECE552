//module ifid(input clk, flush, rst, write, stall_in, input[2:0] ifid_nvz, input[15:0] inst_data, pc, output ifid_flush, stall_out, output [15:0]inst_data_pl, pc_pl);

//wire flush_or_rst;
//assign flush_or_rst = flush | stall_in;
//register_16b pc_reg(.clk(clk), .rst(stall_in |flush ), .write_en(write), .data_in(pc), .data_out(pc_pl));
//register_16b inst_reg(.clk(clk), .rst(stall_in |flush), .write_en(write), .data_in(inst_data), .data_out(inst_data_pl));

//dff flushff(.q(ifid_flush), .d(flush), .wen(write), .clk(clk), .rst(stall_in));
//dff stallff(.q(stall_out), .d(stall_in), .wen(1'b1), .clk(clk), .rst(rst));

//module ifid(input clk, flush, rst, write, input[2:0] ifid_nvz, input[15:0] inst_data, pc, output ifid_flush, output [15:0]inst_data_pl, pc_pl);
module ifid(input clk, flush, rst, write, stall_in, input[2:0] ifid_nvz, input[15:0] inst_data, pc, output ifid_flush, stall_out, output [15:0]inst_data_pl, pc_pl);

wire flush_or_rst;
assign flush_or_rst = flush | rst;
register_16b pc_reg(.clk(clk), .rst(rst |flush ), .write_en(write), .data_in(pc), .data_out(pc_pl));
register_16b inst_reg(.clk(clk), .rst(rst |flush), .write_en(write), .data_in(inst_data), .data_out(inst_data_pl));

dff flushff(.q(ifid_flush), .d(flush), .wen(write), .clk(clk), .rst(rst));
dff stallff(.q(stall_out), .d(stall_in), .wen(write), .clk(clk), .rst(rst));

endmodule

