module dcache(clk, rst_n, address, data_in, enable, mem_wr, write, mem_data_valid, memory_address, data_out, filling_cache, miss_detected);

input clk, rst_n, mem_data_valid, write, enable;
input [15:0] address, data_in;
output [15:0] memory_address, data_out;
output filling_cache, miss_detected;
input mem_wr; // asserted for one clock cycle and passed to memory module

wire miss_detected;
wire [15:0] cache_data_address, memory_address_fsm;
cache_fill_fsm fsm(.clk(clk), .rst_n(rst_n), .miss_address(address & 16'hFFF0), .memory_data_valid(mem_data_valid), .miss_detected(miss_detected), .write_tag_array(write_tag_array),
			.memory_address(memory_address_fsm), .data_address(cache_data_address), .write_data_array(write_data_array), .fsm_busy(filling_cache));

//ouput address for write inst to mem/cache
assign memory_address = (miss_detected) ? memory_address_fsm : address;

// take the address from the PC and decode it
wire [6:0] index_bits;
wire [127:0] BlockEnable;
assign index_bits = (filling_cache) ? cache_data_address[10:4] : address[10:4];
decoder_7_128 block_decoder(.block_address(index_bits), .block(BlockEnable));

// take the address from the PC and choose which word is enabled
wire [2:0] offset_bits;
wire [7:0] WordEnable;
assign offset_bits = (filling_cache) ? cache_data_address[3:1] : address[3:1];
// Cache write: WriteEnable = 1, enable = 1
// Cache read:	WriteEnable = 0, enable = 1
decoder_3_8 word_decoder(.index(offset_bits), .onehot_enable(WordEnable));

//DCACHE: data update writeback
//assign mem_wr =  ~miss_detected; //mem_wr signals memory that it will be written to, send to mem
wire mem_write;
assign mem_write = ~(miss_detected | filling_cache) & mem_wr;
assign cache_wr = miss_detected ? write_data_array : mem_write; //enable cache wr

// cache blocks
wire [15:0] cached_instruction;
DataArray cache_blocks(.clk(clk), .rst(~rst_n), .DataIn(data_in), .Write(cache_wr), .BlockEnable(BlockEnable), .WordEnable(WordEnable), .DataOut(cached_instruction));
assign data_out = (~write_data_array) ? cached_instruction : 16'h0000;

// cache meta
wire [7:0] meta_out, valid_tag;
assign valid_tag = {3'b100, address[15:11]}; // ? is there ever a time when the data in the cache is invalid?
MetaDataArray cache_meta(.clk(clk), .rst(~rst_n), .DataIn(valid_tag), .Write(write_tag_array), .BlockEnable(BlockEnable), .DataOut(meta_out));

// miss detected when the valid bit isn't set or tag bits don't match those for the decoded cache block and word
assign miss_detected = enable & (~meta_out[7] | ~(address[15:11] == meta_out[4:0]));

endmodule
