module  control(input[3:0] opcode, output mem_enable, mem_write);
	
endmodule